
/*
	Christopher Lam
	EE271A
	12/7
	Lab 6
	trees module
	
	This module controls the trees movement, it takes in reset logic from birdwin, outputs 16 bit rows for the led display. 
*/

module trees(clock, reset, start, treein, treein2, treein3, treespass, win, die, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16);

	input logic clock, reset, start, win, die; //single bit logic
	input logic [15:0] treein, treein2, treein3; //16 bit tree logic
	
	output logic [15:0] g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16;//16 bit green rows array
	
	output logic treespass; //output single bit treespass for when all trees have passed the bird
	
	logic [9:0] count; //10 bit logic for counter to slow down logic
	
	enum{S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10, S11, S12, S13, S14, S15, S16, S17, S18, S19, S20, S21, S22, S23, S24, S25} ps, ns; //declare states
	
	//always comb to move trees from one side of the LED array to the other side
	always_comb begin
		case(ps)
			S0: ns = S1;
			S1: ns = S2;
			S2: ns = S3;
			S3: ns = S4;
			S4: ns = S5;
			S5: ns = S6;
			S6: ns = S7;
			S7: ns = S8;
			S8: ns = S9;
			S9: ns = S10;
			S10: ns = S11;
			S11: ns = S12;
			S12: ns = S13;
			S13: ns = S14;
			S14: ns = S15;
			S15: ns = S16;
			S16: ns = S17;
			S17: ns = S18;
			S18: ns = S19;
			S19: ns = S20;
			S20: ns = S21;
			S21: ns = S22;
			S22: ns = S23;
			S23: ns = S24;
			S24: ns = S25;
			S25: ns = S25;
			
		endcase
		
		
		//hard code for different cases, could not figure out how to do this without hard code. 
		case(ps)
		
		S0: begin
			g16 = treein;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S1: begin 
			g16 = 16'b0000000000000000;
			g15 = treein;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S2: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = treein;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S3: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = treein;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S4: begin
			g16 = treein2;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = treein;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S5: begin
			g16 = 16'b0000000000000000;
			g15 = treein2;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = treein;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S6: begin 
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = treein2;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = treein;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S7: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = treein2;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = treein;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S8:begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = treein2;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = treein;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S9: begin
			g16 = treein3;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = treein2;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = treein;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S10: begin
			g16 = 16'b0000000000000000;
			g15 = treein3;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = treein2;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = treein;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S11: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = treein3;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = treein2;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = treein;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S12: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = treein3;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = treein2;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = treein;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S13: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = treein3;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = treein2;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = treein;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S14: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = treein3;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = treein2;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = treein;
		 	g1 = 16'b0000000000000000;
			end
			
		S15: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = treein3;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = treein2;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = treein;
			end
		
		S16: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = treein3;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = treein2;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S17: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = treein3;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = treein2;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S18: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = treein3;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = treein2;
		 	g1 = 16'b0000000000000000;
			end
			
		S19: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = treein3;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = treein2;
			end
			
		S20: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = treein3;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S21: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = treein3;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S22: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = treein3;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		S23: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = treein3;
		 	g1 = 16'b0000000000000000;
			end
			
		S24: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = treein3;
			end
				
		//at this point all trees should have passed the bird
		S25: begin
			g16 = 16'b0000000000000000;
			g15 = 16'b0000000000000000;
			g14 = 16'b0000000000000000;
			g13 = 16'b0000000000000000;
			g12 = 16'b0000000000000000;
		 	g11 = 16'b0000000000000000;
		 	g10 = 16'b0000000000000000;
		 	g9 = 16'b0000000000000000;
		 	g8 = 16'b0000000000000000;
		 	g7 = 16'b0000000000000000;
		 	g6 = 16'b0000000000000000;
		 	g5 = 16'b0000000000000000;
		 	g4 = 16'b0000000000000000;
		 	g3 = 16'b0000000000000000;
		 	g2 = 16'b0000000000000000;
		 	g1 = 16'b0000000000000000;
			end
			
		endcase
	end
			
	//counter to use to slow down logic for this module		
	always_ff @(posedge clock) begin
		if(reset)
			count <= 10'b0000000000;
			
		else if (count == 10'b1111111111)
			count <= 10'b0000000000;
		
		else
			count <= count + 10'b0000000001;
	end	
		
	//reset logic if reset then trees should go back to the beginning side
	always_ff @(posedge clock) begin
		if (reset) begin
			ps <= S0;
			treespass <= 0; //treespass should go back to zero because it goes back to not having passed the bird
		end
		
		else if (win|die) begin //if player wins or dies then reset the trees as well
				ps <= S0;
				treespass <= 0; //same as before
		end
		
		else if (ps == S25) begin //logic to know when the trees have passed the bird, if it makes it to state 25 then it has passed the bird. 
					treespass <= 1;
				end
		
		else if (start) begin //logic to pause the game
			if (count == 10'b1000000000) begin //when count reaches a certain point move to next state, mainly to slow down the logic and actually see it on the display
				ps<=ns;
			
			end
				
		end
		
	end
				
		
		
		
		
		
		
endmodule 

module trees_testbench(); //testbench module for trees

	logic clock, reset, start, treespass, win, die;
	logic [15:0] treein, treein2, treein3;
	
	logic [15:0] g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16;
	
	logic [15:0] out; 
	
	
	trees dut(.clock, .reset, .start, .treein, .treein2, .treein3, .treespass, .win, .die, .g1, .g2, .g3, .g4, .g5, .g6, .g7, .g8, .g9, .g10, .g11, .g12, .g13, .g14, .g15, .g16);
	
	parameter clock_period = 100;
		
			initial begin
				clock <= 0;
				forever #(clock_period /2) clock <= ~clock; //every 100/2 period flip the bit of the clock set by DE1_SoC
					
			end 
		
			initial begin //manually set inputs for pattern
		
			reset <= 1; 																@(posedge clock);//reset once
			reset <= 0; start <= 1; treein <= 16'b1111110001111111; 		@(posedge clock);//set reset to 0, and unpause game
																							@(posedge clock);
																							@(posedge clock);//tree should be moving
																							@(posedge clock);
											treein2 <= 16'b1111110001111111;		@(posedge clock);//second tree
																							@(posedge clock);
																							@(posedge clock);
																								@(posedge clock);
											treein3 <= 16'b1111110001111111;		@(posedge clock); //third tree
																								@(posedge clock);
																							@(posedge clock);
																								@(posedge clock);
																							@(posedge clock);
																							@(posedge clock);
																								@(posedge clock);	
																								@(posedge clock);
																								@(posedge clock);	
																							@(posedge clock);
																							@(posedge clock);
			$stop; //end simulation							
							
		end 
		
endmodule		
			
			